* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d0 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nch_lvt_mac_CDNS_579155404420 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch_lvt L=6e-08 W=2e-07 $X=0 $Y=0 $D=46
.ENDS
***************************************
.SUBCKT nch_lvt_mac_CDNS_579155404421 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch_lvt L=6e-08 W=2e-07 $X=0 $Y=0 $D=46
.ENDS
***************************************
.SUBCKT currentmirror_single_n S0 D G
** N=3 EP=3 IP=8 FDC=2
X0 S0 D G S0 nch_lvt_mac_CDNS_579155404420 $T=100 340 0 0 $X=-295 $Y=0
X1 D S0 G S0 nch_lvt_mac_CDNS_579155404421 $T=360 340 0 0 $X=-35 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3
** N=3 EP=3 IP=6 FDC=4
X0 1 3 2 currentmirror_single_n $T=0 0 0 0 $X=-295 $Y=-90
X1 1 3 2 currentmirror_single_n $T=520 0 0 0 $X=225 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3
** N=3 EP=3 IP=6 FDC=8
X0 1 2 3 ICV_1 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_1 $T=1040 0 0 0 $X=745 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3
** N=3 EP=3 IP=6 FDC=16
X0 1 2 3 ICV_2 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_2 $T=2080 0 0 0 $X=1785 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3
** N=3 EP=3 IP=6 FDC=32
X0 1 2 3 ICV_3 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_3 $T=4160 0 0 0 $X=3865 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3
** N=3 EP=3 IP=6 FDC=64
X0 1 2 3 ICV_4 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_4 $T=8320 0 0 0 $X=8025 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3
** N=3 EP=3 IP=6 FDC=128
X0 1 2 3 ICV_5 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_5 $T=16640 0 0 0 $X=16345 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3
** N=3 EP=3 IP=6 FDC=256
X0 1 2 3 ICV_6 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 ICV_6 $T=33280 0 0 0 $X=32985 $Y=-90
.ENDS
***************************************
.SUBCKT diffpair_two_finger_n S0 D S1 G 5
** N=5 EP=5 IP=8 FDC=2
X0 S0 D G 5 nch_lvt_mac_CDNS_579155404420 $T=100 140 0 0 $X=-295 $Y=-200
X1 D S1 G 5 nch_lvt_mac_CDNS_579155404421 $T=360 140 0 0 $X=-35 $Y=-200
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4
** N=4 EP=4 IP=10 FDC=4
X0 1 3 1 2 4 diffpair_two_finger_n $T=0 0 0 0 $X=-295 $Y=-200
X1 1 3 1 2 4 diffpair_two_finger_n $T=520 0 0 0 $X=225 $Y=-200
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=8
X0 1 3 2 ICV_1 $T=0 0 0 0 $X=-295 $Y=-90
X1 2 4 5 1 ICV_8 $T=0 2030 0 0 $X=-295 $Y=1830
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=16
X0 1 2 3 4 5 ICV_9 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_9 $T=1040 0 0 0 $X=745 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=32
X0 1 2 3 4 5 ICV_10 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_10 $T=2080 0 0 0 $X=1785 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=64
X0 1 2 3 4 5 ICV_11 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_11 $T=4160 0 0 0 $X=3865 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=128
X0 1 2 3 4 5 ICV_12 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_12 $T=8320 0 0 0 $X=8025 $Y=-90
.ENDS
***************************************
.SUBCKT activeload_two_finger_p S0 D S1 G 6
** N=6 EP=5 IP=0 FDC=2
M0 D G S0 6 pch_lvt L=6e-08 W=2e-07 $X=100 $Y=240 $D=118
M1 S1 G D 6 pch_lvt L=6e-08 W=2e-07 $X=360 $Y=240 $D=118
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3
** N=4 EP=3 IP=12 FDC=4
X0 2 3 2 1 2 activeload_two_finger_p $T=0 0 0 0 $X=-390 $Y=-380
X1 2 3 2 1 2 activeload_two_finger_p $T=520 0 0 0 $X=130 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3
** N=4 EP=3 IP=8 FDC=8
X0 1 2 3 ICV_14 $T=0 0 0 0 $X=-390 $Y=-380
X1 1 2 3 ICV_14 $T=1040 0 0 0 $X=650 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7
** N=7 EP=7 IP=9 FDC=24
X0 1 2 3 4 7 ICV_10 $T=0 0 0 0 $X=-295 $Y=-90
X1 5 6 7 ICV_15 $T=0 4060 0 0 $X=-390 $Y=3680
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7
** N=7 EP=7 IP=14 FDC=48
X0 1 2 3 4 5 6 7 ICV_16 $T=0 0 0 0 $X=-390 $Y=-90
X1 1 2 3 4 5 6 7 ICV_16 $T=2080 0 0 0 $X=1690 $Y=-90
.ENDS
***************************************
.SUBCKT currentmirror_ref_n S0 D
** N=2 EP=2 IP=8 FDC=2
X0 S0 D D S0 nch_lvt_mac_CDNS_579155404420 $T=100 340 0 0 $X=-295 $Y=0
X1 D S0 D S0 nch_lvt_mac_CDNS_579155404421 $T=360 340 0 0 $X=-35 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT ICV_18 1 2
** N=2 EP=2 IP=4 FDC=4
X0 1 2 currentmirror_ref_n $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 currentmirror_ref_n $T=520 0 0 0 $X=225 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 ICV_18 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_18 $T=1040 0 0 0 $X=745 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_20 1 2
** N=2 EP=2 IP=4 FDC=16
X0 1 2 ICV_19 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_19 $T=2080 0 0 0 $X=1785 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_21 1 2
** N=2 EP=2 IP=4 FDC=32
X0 1 2 ICV_20 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_20 $T=4160 0 0 0 $X=3865 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_22 1 2
** N=2 EP=2 IP=4 FDC=64
X0 1 2 ICV_21 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_21 $T=8320 0 0 0 $X=8025 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=4 FDC=128
X0 1 2 ICV_22 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_22 $T=16640 0 0 0 $X=16345 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_24 1 2
** N=2 EP=2 IP=4 FDC=256
X0 1 2 ICV_23 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 ICV_23 $T=33280 0 0 0 $X=32985 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=8
X0 1 3 5 2 ICV_8 $T=0 2030 0 0 $X=-295 $Y=1830
X1 2 4 ICV_18 $T=0 0 0 0 $X=-295 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=16
X0 2 1 4 3 5 ICV_25 $T=0 0 0 0 $X=-295 $Y=-90
X1 2 1 4 3 5 ICV_25 $T=1040 0 0 0 $X=745 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=32
X0 1 2 3 4 5 ICV_26 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_26 $T=2080 0 0 0 $X=1785 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=64
X0 1 2 3 4 5 ICV_27 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_27 $T=4160 0 0 0 $X=3865 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5
** N=5 EP=5 IP=10 FDC=128
X0 1 2 3 4 5 ICV_28 $T=0 0 0 0 $X=-295 $Y=-90
X1 1 2 3 4 5 ICV_28 $T=8320 0 0 0 $X=8025 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7
** N=7 EP=7 IP=9 FDC=24
X0 3 4 7 ICV_15 $T=0 4060 0 0 $X=-390 $Y=3680
X1 1 2 5 6 7 ICV_26 $T=0 0 0 0 $X=-295 $Y=-90
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7
** N=7 EP=7 IP=14 FDC=48
X0 1 2 5 6 3 4 7 ICV_30 $T=0 0 0 0 $X=-390 $Y=-90
X1 1 2 5 6 3 4 7 ICV_30 $T=2080 0 0 0 $X=1690 $Y=-90
.ENDS
***************************************
.SUBCKT DIFFAMP_lch_60n VSS VDD inm vbias inp idc outp outm
** N=9 EP=8 IP=223 FDC=5868
X0 VSS idc 3 ICV_3 $T=1181960 0 0 0 $X=1181665 $Y=-90
X1 VSS idc 3 ICV_4 $T=1173640 0 0 0 $X=1173345 $Y=-90
X2 VSS idc 3 ICV_6 $T=1140360 0 0 0 $X=1140065 $Y=-90
X3 VSS idc 3 ICV_7 $T=741000 0 0 0 $X=740705 $Y=-90
X4 VSS idc 3 ICV_7 $T=807560 0 0 0 $X=807265 $Y=-90
X5 VSS idc 3 ICV_7 $T=874120 0 0 0 $X=873825 $Y=-90
X6 VSS idc 3 ICV_7 $T=940680 0 0 0 $X=940385 $Y=-90
X7 VSS idc 3 ICV_7 $T=1007240 0 0 0 $X=1006945 $Y=-90
X8 VSS idc 3 ICV_7 $T=1073800 0 0 0 $X=1073505 $Y=-90
X9 3 outp 3 inm VSS diffpair_two_finger_n $T=147680 2030 0 0 $X=147385 $Y=1830
X10 3 outm 3 inp VSS diffpair_two_finger_n $T=741000 2030 0 0 $X=740705 $Y=1830
X11 VSS 3 idc inp outm ICV_10 $T=738920 0 0 0 $X=738625 $Y=-90
X12 VSS 3 idc inp outm ICV_12 $T=730600 0 0 0 $X=730305 $Y=-90
X13 VSS 3 idc inp outm ICV_13 $T=614120 0 0 0 $X=613825 $Y=-90
X14 VSS 3 idc inp outm ICV_13 $T=630760 0 0 0 $X=630465 $Y=-90
X15 VSS 3 idc inp outm ICV_13 $T=647400 0 0 0 $X=647105 $Y=-90
X16 VSS 3 idc inp outm ICV_13 $T=664040 0 0 0 $X=663745 $Y=-90
X17 VSS 3 idc inp outm ICV_13 $T=680680 0 0 0 $X=680385 $Y=-90
X18 VSS 3 idc inp outm ICV_13 $T=697320 0 0 0 $X=697025 $Y=-90
X19 VSS 3 idc inp outm ICV_13 $T=713960 0 0 0 $X=713665 $Y=-90
X20 vbias VDD outp ICV_14 $T=20800 4060 0 0 $X=20410 $Y=3680
X21 vbias VDD outm ICV_14 $T=614120 4060 0 0 $X=613730 $Y=3680
X22 VSS 3 idc inp vbias VDD outm ICV_17 $T=593320 0 0 0 $X=592930 $Y=-90
X23 VSS 3 idc inp vbias VDD outm ICV_17 $T=597480 0 0 0 $X=597090 $Y=-90
X24 VSS 3 idc inp vbias VDD outm ICV_17 $T=601640 0 0 0 $X=601250 $Y=-90
X25 VSS 3 idc inp vbias VDD outm ICV_17 $T=605800 0 0 0 $X=605410 $Y=-90
X26 VSS 3 idc inp vbias VDD outm ICV_17 $T=609960 0 0 0 $X=609570 $Y=-90
X27 VSS idc ICV_20 $T=588640 0 0 0 $X=588345 $Y=-90
X28 VSS idc ICV_21 $T=580320 0 0 0 $X=580025 $Y=-90
X29 VSS idc ICV_23 $T=547040 0 0 0 $X=546745 $Y=-90
X30 VSS idc ICV_24 $T=147680 0 0 0 $X=147385 $Y=-90
X31 VSS idc ICV_24 $T=214240 0 0 0 $X=213945 $Y=-90
X32 VSS idc ICV_24 $T=280800 0 0 0 $X=280505 $Y=-90
X33 VSS idc ICV_24 $T=347360 0 0 0 $X=347065 $Y=-90
X34 VSS idc ICV_24 $T=413920 0 0 0 $X=413625 $Y=-90
X35 VSS idc ICV_24 $T=480480 0 0 0 $X=480185 $Y=-90
X36 VSS 3 idc inm outp ICV_26 $T=145600 0 0 0 $X=145305 $Y=-90
X37 VSS 3 idc inm outp ICV_28 $T=137280 0 0 0 $X=136985 $Y=-90
X38 VSS 3 idc inm outp ICV_29 $T=20800 0 0 0 $X=20505 $Y=-90
X39 VSS 3 idc inm outp ICV_29 $T=37440 0 0 0 $X=37145 $Y=-90
X40 VSS 3 idc inm outp ICV_29 $T=54080 0 0 0 $X=53785 $Y=-90
X41 VSS 3 idc inm outp ICV_29 $T=70720 0 0 0 $X=70425 $Y=-90
X42 VSS 3 idc inm outp ICV_29 $T=87360 0 0 0 $X=87065 $Y=-90
X43 VSS 3 idc inm outp ICV_29 $T=104000 0 0 0 $X=103705 $Y=-90
X44 VSS 3 idc inm outp ICV_29 $T=120640 0 0 0 $X=120345 $Y=-90
X45 VSS 3 idc inm vbias VDD outp ICV_31 $T=0 0 0 0 $X=-390 $Y=-90
X46 VSS 3 idc inm vbias VDD outp ICV_31 $T=4160 0 0 0 $X=3770 $Y=-90
X47 VSS 3 idc inm vbias VDD outp ICV_31 $T=8320 0 0 0 $X=7930 $Y=-90
X48 VSS 3 idc inm vbias VDD outp ICV_31 $T=12480 0 0 0 $X=12090 $Y=-90
X49 VSS 3 idc inm vbias VDD outp ICV_31 $T=16640 0 0 0 $X=16250 $Y=-90
.ENDS
***************************************
