* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d0 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nch_lvt_mac_CDNS_583293706990 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch_lvt L=6e-08 W=2e-07 $X=0 $Y=0 $D=46
.ENDS
***************************************
.SUBCKT nch_lvt_mac_CDNS_583293706991 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch_lvt L=6e-08 W=2e-07 $X=0 $Y=0 $D=46
.ENDS
***************************************
.SUBCKT currentmirror_single_n D G S0
** N=3 EP=3 IP=8 FDC=2
X0 S0 D G S0 nch_lvt_mac_CDNS_583293706990 $T=100 340 0 0 $X=-295 $Y=0
X1 D S0 G S0 nch_lvt_mac_CDNS_583293706991 $T=360 340 0 0 $X=-35 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT diffpair_two_finger_n D G S0 S1 5
** N=5 EP=5 IP=8 FDC=2
X0 S0 D G 5 nch_lvt_mac_CDNS_583293706990 $T=100 140 0 0 $X=-295 $Y=-200
X1 D S1 G 5 nch_lvt_mac_CDNS_583293706991 $T=360 140 0 0 $X=-35 $Y=-200
.ENDS
***************************************
.SUBCKT activeload_two_finger_p S0 D S1 G 6
** N=6 EP=5 IP=0 FDC=2
M0 D G S0 6 pch_lvt L=6e-08 W=2e-07 $X=100 $Y=240 $D=118
M1 S1 G D 6 pch_lvt L=6e-08 W=2e-07 $X=360 $Y=240 $D=118
.ENDS
***************************************
.SUBCKT currentmirror_ref_n D S0
** N=2 EP=2 IP=8 FDC=2
X0 S0 D D S0 nch_lvt_mac_CDNS_583293706990 $T=100 340 0 0 $X=-295 $Y=0
X1 D S0 D S0 nch_lvt_mac_CDNS_583293706991 $T=360 340 0 0 $X=-35 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT DIFFAMP_lch_60n VSS VDD inm vbias inp idc outp outm
** N=9 EP=8 IP=84 FDC=48
X0 7 idc VSS currentmirror_single_n $T=4680 0 0 0 $X=4385 $Y=-90
X1 7 idc VSS currentmirror_single_n $T=5200 0 0 0 $X=4905 $Y=-90
X2 7 idc VSS currentmirror_single_n $T=5720 0 0 0 $X=5425 $Y=-90
X3 7 idc VSS currentmirror_single_n $T=6240 0 0 0 $X=5945 $Y=-90
X4 7 idc VSS currentmirror_single_n $T=6760 0 0 0 $X=6465 $Y=-90
X5 7 idc VSS currentmirror_single_n $T=7280 0 0 0 $X=6985 $Y=-90
X6 7 idc VSS currentmirror_single_n $T=7800 0 0 0 $X=7505 $Y=-90
X7 7 idc VSS currentmirror_single_n $T=8320 0 0 0 $X=8025 $Y=-90
X8 outp inm 7 7 VSS diffpair_two_finger_n $T=0 2030 0 0 $X=-295 $Y=1830
X9 outp inm 7 7 VSS diffpair_two_finger_n $T=520 2030 0 0 $X=225 $Y=1830
X10 outm inp 7 7 VSS diffpair_two_finger_n $T=4680 2030 0 0 $X=4385 $Y=1830
X11 outm inp 7 7 VSS diffpair_two_finger_n $T=5200 2030 0 0 $X=4905 $Y=1830
X12 VDD outp VDD vbias VDD activeload_two_finger_p $T=0 4060 0 0 $X=-390 $Y=3680
X13 VDD outp VDD vbias VDD activeload_two_finger_p $T=520 4060 0 0 $X=130 $Y=3680
X14 VDD outm VDD vbias VDD activeload_two_finger_p $T=4680 4060 0 0 $X=4290 $Y=3680
X15 VDD outm VDD vbias VDD activeload_two_finger_p $T=5200 4060 0 0 $X=4810 $Y=3680
X16 idc VSS currentmirror_ref_n $T=0 0 0 0 $X=-295 $Y=-90
X17 idc VSS currentmirror_ref_n $T=520 0 0 0 $X=225 $Y=-90
X18 idc VSS currentmirror_ref_n $T=1040 0 0 0 $X=745 $Y=-90
X19 idc VSS currentmirror_ref_n $T=1560 0 0 0 $X=1265 $Y=-90
X20 idc VSS currentmirror_ref_n $T=2080 0 0 0 $X=1785 $Y=-90
X21 idc VSS currentmirror_ref_n $T=2600 0 0 0 $X=2305 $Y=-90
X22 idc VSS currentmirror_ref_n $T=3120 0 0 0 $X=2825 $Y=-90
X23 idc VSS currentmirror_ref_n $T=3640 0 0 0 $X=3345 $Y=-90
.ENDS
***************************************
